module im(
input [31:0]address,
input en,
output [31:0]inst_out);

reg[31:0] inst_mem[31:0];

initial
begin
//R TYPE
inst_mem[0]=32'b0;
inst_mem[1]=32'b0000001_00001_00000_000_10101_0110011;//MUL
inst_mem[2]=32'b0000001_00010_00000_001_10101_0110011;//MULH
inst_mem[3]=32'b0000001_00011_00000_010_10101_0110011;//MULHSU
inst_mem[4]=32'b0000001_00100_00000_011_10101_0110011;//MULHU
inst_mem[5]=32'b0000001_00101_00000_100_10101_0110011;//DIV
inst_mem[6]=32'b0000001_00110_00000_101_10101_0110011;//DIVU
inst_mem[7]=32'b0000001_00111_00000_110_10101_0110011;//REM
inst_mem[8]=32'b0000001_01000_00000_111_10101_0110011;//REMU
inst_mem[9]=32'b0000000_00010_00001_000_00101_0110011;//ADD
inst_mem[10]=32'b0100000_00100_00011_000_00110_0110011;//SUB
inst_mem[11]=32'b0000000_00110_00101_111_00111_0110011;//AND
inst_mem[12]=32'b0000000_00010_00001_110_01000_0110011;//OR
inst_mem[13]=32'b0000000_00011_00010_100_01001_0110011;//XOR
inst_mem[14]=32'b0000000_00010_00001_001_01010_0110011;//SLL
inst_mem[15]=32'b0000000_00010_00001_101_01011_0110011;//SRL
inst_mem[16]=32'b0100000_00010_00001_101_01100_0110011;//SRA
inst_mem[17]=32'b0000000_00010_00001_010_01101_0110011;//SLT


//I TYPE
inst_mem[18]=32'b000000000011_00001_000_00001_0010011;//addi
inst_mem[19]=32'b000000001000_00010_111_00010_0010011;//andi
inst_mem[20]=32'b000000000001_00011_110_00011_0010011;//ori
inst_mem[21]=32'b000000000010_00100_100_00100_0010011;//xori
inst_mem[22]=32'b000000000101_00010_010_01001_0010011;//SLTI
inst_mem[23]=32'b000000000101_00010_011_01001_0010011;//SLTIU
inst_mem[24]=32'b000000000010_00001_001_01011_0010011;//SLLI
inst_mem[25]=32'b000000000011_00001_101_01100_0010011;//SRLI
inst_mem[26]=32'b010000000100_00001_101_01101_0010011;//SRAI


//S TYPE
inst_mem[27]=32'b0000000_00110_00010_010_01100_0100011;//SW
inst_mem[28]=32'b0000000_00111_00011_001_00100_0100011;//SH
inst_mem[29]=32'b0000000_01000_00100_000_00000_0100011;//SB


//U TYPE
inst_mem[30]=32'b000010010001101000101_01010_0110111;//LUI
inst_mem[31]=32'b000010010001101000101_01010_0010111;//AUIPC



end


assign inst_out = (en) ? inst_mem[address]:32'b0;

endmodule 

